module top_module( input in, output out );
assign out=~in;
endmodule

//this module is used to define just working of a NOT gate or an Inverter
